module FSM_SAW (
    
);
    
endmodule